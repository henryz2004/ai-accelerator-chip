module packet_io #(
	parameter fifo_len=4,
	parameter max_data_bytes=8
)
(

);

endmodule 